library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

entity cos is
    port 
    (
        u,x : in unsigned(2 downto 0);  
        c : out sfixed(1 downto -16) --c is cos in signed fixed point
    ) ;
end cos;

architecture arch of cos is

    signal  ux: UNSIGNED(5 downto 0);
begin
    ux <= u&x;
    with ux select
    c <=
    "010000000000000000" when "000000",
    "010000000000000000" when "000001",
    "010000000000000000" when "000010",
    "010000000000000000" when "000011",
    "010000000000000000" when "000100",
    "010000000000000000" when "000101",
    "010000000000000000" when "000110",
    "010000000000000000" when "000111",
    "110000010011000011" when "001000",
    "110010101101000100" when "001001",
    "110111000110101001" when "001010",
    "111100111000010101" when "001011",
    "000011000111101011" when "001100",
    "001000111001010111" when "001101",
    "001101010010111100" when "001110",
    "001111101100111101" when "001111",
    "001110110011110110" when "010000",
    "000111010001111010" when "010001",
    "111000101110000110" when "010010",
    "110001001100001010" when "010011",
    "110001001100001010" when "010100",
    "111000101110000110" when "010101",
    "000111010001111010" when "010110",
    "001110110011110110" when "010111",
    "110010101101000100" when "011000",
    "000011000111101011" when "011001",
    "001111101100111101" when "011010",
    "001000111001010111" when "011011",
    "110111000110101001" when "011100",
    "110000010011000011" when "011101",
    "111100111000010101" when "011110",
    "001101010010111100" when "011111",
    "001011010011111101" when "100000",
    "110100101100000011" when "100001",
    "110100101100000011" when "100010",
    "001011010011111101" when "100011",
    "001011010011111101" when "100100",
    "110100101100000011" when "100101",
    "110100101100000011" when "100110",
    "001011010011111101" when "100111",
    "110111000110101001" when "101000",
    "001111101100111101" when "101001",
    "111100111000010101" when "101010",
    "110010101101000100" when "101011",
    "001101010010111100" when "101100",
    "000011000111101011" when "101101",
    "110000010011000011" when "101110",
    "001000111001010111" when "101111",
    "000111010001111010" when "110000",
    "110001001100001010" when "110001",
    "001110110011110110" when "110010",
    "111000101110000110" when "110011",
    "111000101110000110" when "110100",
    "001110110011110110" when "110101",
    "110001001100001010" when "110110",
    "000111010001111010" when "110111",
    "111100111000010101" when "111000",
    "001000111001010111" when "111001",
    "110010101101000100" when "111010",
    "001111101100111101" when "111011",
    "110000010011000011" when "111100",
    "001101010010111100" when "111101",
    "110111000110101001" when "111110",
    "000011000111101011" when "111111";

end arch ; -- arch