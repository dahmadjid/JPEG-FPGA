library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;



package jpeg_pkg is 
    
    type image_row_t is array (0 to 7) of unsigned(7 downto 0);
    type image_block_t is array (0 to 7) of image_row_t; --8 by 8 block of image
    type qz_row_t is array (0 to 7) of ufixed(16 downto 0);
    type qz_table_t is array (0 to 7) of qz_row_t;
    type dct_coeff_row_t is array(0 to 7) of sfixed(10 downto 0);
    type dct_coeff_block_t is array(0 to 7) of dct_coeff_row_t; --8 by 8 dct coeff array
    -- type dct_coeff_yx_row_t is array(0 to 7) of sfixed(13 downto -32);
    -- type dct_coeff_yx_mat_t is array(0 to 7) of dct_coeff_yx_row_t;
    type cos_row_t is array(0 to 7) of sfixed(1 downto -16);
    type cos_mat_t is array(0 to 7) of cos_row_t;
    -- constant luminance_qz: image_block_t := 
    -- ("00010000","00001011","00001010","00010000","00011000","00101000","00110011","00111101"),
    -- ("00001100","00001100","00001110","00010011","00011010","00111010","00111100","00110111"),
    -- ("00001110","00001101","00010000","00011000","00101000","00111001","01000101","00111000"),
    -- ("00001110","00010001","00010110","00011101","00110011","01010111","01010000","00111110"),
    -- ("00010010","00010110","00100101","00111000","01000100","01101101","01100111","01001101"),
    -- ("00011000","00100011","00110111","01000000","01010001","01101000","01110001","01011100"),
    -- ("00110001","01000000","01001110","01010111","01100111","01111001","01111000","01100101"),
    -- ("01001000","01011100","01011111","01100010","01110000","01100100","01100111","01100011");
    
    -- constant chrominance_qz: image_block_t := 
    -- ("00010001","00010010","00011000","00101111","01100011","01100011","01100011","01100011"),
    -- ("00010010","00010101","00011010","01000010","01100011","01100011","01100011","01100011"),
    -- ("00011000","00011010","00111000","01100011","01100011","01100011","01100011","01100011"),
    -- ("00101111","01000010","01100011","01100011","01100011","01100011","01100011","01100011"),
    -- ("01100011","01100011","01100011","01100011","01100011","01100011","01100011","01100011"),
    -- ("01100011","01100011","01100011","01100011","01100011","01100011","01100011","01100011"),
    -- ("01100011","01100011","01100011","01100011","01100011","01100011","01100011","01100011"),
    -- ("01100011","01100011","01100011","01100011","01100011","01100011","01100011","01100011");
    
    -- constant luminance_qz_shift: qz_table_t := 
    -- ("0000111111111111","0001011101000101","0001100110011001","0000111111111111","0000101010101010","0000011001100110","0000010100000101","0000010000110010"),
    -- ("0001010101010101","0001010101010101","0001001001001001","0000110101111001","0000100111011000","0000010001101001","0000010001000100","0000010010100111"),
    -- ("0001001001001001","0001001110110001","0000111111111111","0000101010101010","0000011001100110","0000010001111101","0000001110110101","0000010010010010"),
    -- ("0001001001001001","0000111100001111","0000101110100010","0000100011010011","0000010100000101","0000001011110001","0000001100110011","0000010000100001"),
    -- ("0000111000111000","0000101110100010","0000011011101011","0000010010010010","0000001111000011","0000001001011001","0000001001111100","0000001101010011"),
    -- ("0000101010101010","0000011101010000","0000010010100111","0000001111111111","0000001100101001","0000001001110110","0000001001000011","0000001011001000"),
    -- ("0000010100111001","0000001111111111","0000001101001000","0000001011110001","0000001001111100","0000001000011101","0000001000100010","0000001010001000"),
    -- ("0000001110001110","0000001011001000","0000001010110001","0000001010011100","0000001001001001","0000001010001111","0000001001111100","0000001010010101");
    
    -- constant chrominance_qz_shift: qz_table_t := 
    -- ("0000111100001111","0000111000111000","0000101010101010","0000010101110010","0000001010010101","0000001010010101","0000001010010101","0000001010010101"),
    -- ("0000111000111000","0000110000110000","0000100111011000","0000001111100000","0000001010010101","0000001010010101","0000001010010101","0000001010010101"),
    -- ("0000101010101010","0000100111011000","0000010010010010","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101"),
    -- ("0000010101110010","0000001111100000","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101"),
    -- ("0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101"),
    -- ("0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101"),
    -- ("0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101"),
    -- ("0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101","0000001010010101");
    
    component cos is   
        port 
        (
        u,x : in unsigned(2 downto 0);   
        c : out sfixed(1 downto -16)       --c is cos in signed fixed point
        );
    end component;
    component constant_v is  
        port (
        u,x : in unsigned(2 downto 0);
        const : out sfixed(1 downto -16)
        ) ;
    end component;
    component dct is
        port (
            u,v : in unsigned(2 downto 0);
            img_block : in image_block_t;
            dct_coeff : out sfixed(10 downto 0)
          ) ;
    end component;
    component mini_length is
        port 
        (
            dct_coeff : in sfixed(10 downto 0);  
            huff_value : out sfixed(10 downto 0);
            length : out unsigned(3 downto 0) --number between 0 and 11
        ) ;
    end component;
    
    component y_quantizer is
    port (
      dct_coeff_block : in dct_coeff_block_t;
      dct_coeff_qz : out dct_coeff_block_t
    ) ;
    end component;

    component c_quantizer is
    port (
      dct_coeff_block : in dct_coeff_block_t;
      dct_coeff_qz : out dct_coeff_block_t
    ) ;
    end component;
    

end package;