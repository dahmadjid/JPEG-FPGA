library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
-- TESTED IN FPGA. WORKS GOOD
entity cos is
    port 
    (
        u,x : in unsigned(2 downto 0);  
        c : out sfixed(1 downto -20) --c is cos in signed fixed point
    ) ;
end cos;

architecture arch of cos is

    signal  ux: UNSIGNED(5 downto 0);
begin
    ux <= u&x;
    with ux select
    c <= 
    "0100000000000000000000" when "000000",
    "0100000000000000000000" when "000001",
    "0100000000000000000000" when "000010",
    "0100000000000000000000" when "000011",
    "0100000000000000000000" when "000100",
    "0100000000000000000000" when "000101",
    "0100000000000000000000" when "000110",
    "0100000000000000000000" when "000111",
    "0011111011000101001011" when "001000",
    "0011010100110110110011" when "001001",
    "0010001110001110011101" when "001010",
    "0000110001111100010111" when "001011",
    "1111001110000011101001" when "001100",
    "1101110001110001100011" when "001101",
    "1100101011001001001101" when "001110",
    "1100000100111010110101" when "001111",
    "0011101100100000110101" when "010000",
    "0001100001111101111000" when "010001",
    "1110011110000010001000" when "010010",
    "1100010011011111001011" when "010011",
    "1100010011011111001011" when "010100",
    "1110011110000010001000" when "010101",
    "0001100001111101111000" when "010110",
    "0011101100100000110101" when "010111",
    "0011010100110110110011" when "011000",
    "1111001110000011101001" when "011001",
    "1100000100111010110101" when "011010",
    "1101110001110001100011" when "011011",
    "0010001110001110011101" when "011100",
    "0011111011000101001011" when "011101",
    "0000110001111100010111" when "011110",
    "1100101011001001001101" when "011111",
    "0010110101000001001111" when "100000",
    "1101001010111110110001" when "100001",
    "1101001010111110110001" when "100010",
    "0010110101000001001111" when "100011",
    "0010110101000001001111" when "100100",
    "1101001010111110110001" when "100101",
    "1101001010111110110001" when "100110",
    "0010110101000001001111" when "100111",
    "0010001110001110011101" when "101000",
    "1100000100111010110101" when "101001",
    "0000110001111100010111" when "101010",
    "0011010100110110110011" when "101011",
    "1100101011001001001101" when "101100",
    "1111001110000011101001" when "101101",
    "0011111011000101001011" when "101110",
    "1101110001110001100011" when "101111",
    "0001100001111101111000" when "110000",
    "1100010011011111001011" when "110001",
    "0011101100100000110101" when "110010",
    "1110011110000010001000" when "110011",
    "1110011110000010001000" when "110100",
    "0011101100100000110101" when "110101",
    "1100010011011111001011" when "110110",
    "0001100001111101111000" when "110111",
    "0000110001111100010111" when "111000",
    "1101110001110001100011" when "111001",
    "0011010100110110110011" when "111010",
    "1100000100111010110101" when "111011",
    "0011111011000101001011" when "111100",
    "1100101011001001001101" when "111101",
    "0010001110001110011101" when "111110",
    "1111001110000011101001" when "111111";
    
end arch ; -- arch