library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity bram is
  port (
    clock : in std_logic;
    address : in std_logic_vector();


  ) ;
end bram;